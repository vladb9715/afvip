// -----------------------------------------------------------------------------
// Module name: afvip_apb_pkg
// HDL        : System Verilog
// Author     : Vlad Botezatu
// Description: Keep all of the reset components in an organized fashion.
// Date       : 25 July, 2023
// -----------------------------------------------------------------------------
package afvip_rst_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    `include "afvip_rst_item.svh"
    `include "afvip_rst_sequencer.svh"
    `include "afvip_rst_driver.svh"
    `include "afvip_rst_monitor.svh"
    `include "afvip_rst_agent.svh"
    `include "afvip_rst_sequence.svh"
endpackage : afvip_rst_pkg